LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

entity ps2_mouse is
	port
	(
		CLOCK_50		: 		in			STD_LOGIC;											
		reset 		:		in			STD_LOGIC;				
		PS2_DAT 		:		inout		STD_LOGIC;	--	PS2 Data
		PS2_CLK		:		inout		STD_LOGIC;	--	PS2 Clock
		data_mouse	: 		out 		STD_LOGIC_VECTOR (15 downto 0);
		Click			: 		out		STD_LOGIC
	);
end entity;

architecture struct of ps2_mouse is
	
	component mouse_ctrl
		generic(
			clkfreq : integer
		);
		port(
			ps2_data		:	inout	std_logic;
			ps2_clk		:	inout	std_logic;
			clk			:	in 	std_logic;
			en				:	in 	std_logic;
			resetn		:	in 	std_logic;
			newdata		:	out	std_logic;
			bt_on			:	out	std_logic_vector(2 downto 0);
			ox, oy		:	out 	std_logic;
			dx, dy		:	out	std_logic_vector(8 downto 0);
			wheel			: 	out	std_logic_vector(3 downto 0)
		);
	end component;
	
	signal signewdata, resetn : std_logic;
	signal dx, dy : std_logic_vector(8 downto 0);
	signal x, y 	: std_logic_vector(7 downto 0);
	signal data : std_logic_vector(15 downto 0);
	signal botoes : std_logic_vector(2 downto 0);
	signal overflow_x, overflow_y : std_logic;
	signal wheel : std_logic_vector(3 downto 0);
	
	constant SENSIBILITY : integer := 8; -- Rise to decrease sensibility
	
begin 
	resetn <= reset;
	
	mousectrl : mouse_ctrl generic map (50000) port map(
				PS2_DAT,
				PS2_CLK, 
				CLOCK_50,
				'1', 
				reset,
				signewdata, 
				botoes(2 downto 0),
				overflow_x,
				overflow_y,
				dx,
				dy, 
				wheel
	);
	
	-- Read new mouse data	
	process(signewdata, resetn)
		variable xacc, yacc : integer range -10000 to 10000;
	begin
		if(rising_edge(signewdata)) then			
			x <= std_logic_vector(to_signed(to_integer(signed(x)) + ((xacc + to_integer(signed(dx))) / SENSIBILITY), 8));
			y <= std_logic_vector(to_signed(to_integer(signed(y)) + ((yacc + to_integer(signed(dy))) / SENSIBILITY), 8));
			xacc := ((xacc + to_integer(signed(dx))) rem SENSIBILITY);
			yacc := ((yacc + to_integer(signed(dy))) rem SENSIBILITY);					
		end if;
		if resetn = '0' then
			xacc := 0;
			yacc := 0;
			x <= (others => '0');
			y <= (others => '0');
		end if;
	end process;

	data(3  downto  0) <= y(3 downto 0);
	data(7  downto  4) <= y(7 downto 4);
	data(11 downto  8) <= x(3 downto 0);
	data(15 downto 12) <= x(7 downto 4);
	
	data_mouse <= data;
	Click <= botoes(0);

end struct;